
`define c_IIR_NBITS		40
`define c_NUM_REGS		10
`define c_CMD_NBITS  	8
`define c_BUF_NBITS 		48
`define c_ACCUM_NBITS 	72
