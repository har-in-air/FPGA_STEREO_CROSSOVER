
`define c_CMD_NBITS  		8
`define c_COEFF_NBITS		40
`define c_COEFF_FBITS		36
`define c_NCOEFFS				20
`define c_DATA_NBITS			24
`define c_BUF_NBITS 			48
`define c_MULT_NBITS 		64
`define c_ACCUM_NBITS 		72
